library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Decoder is
     Generic( NUMBITS: integer := 32 );
     Port ( clk : in std_logic;
            rst : in std_logic;
            read_in : in std_logic;
            input : in std_logic_vector( 4 downto 0 );
            output : out std_logic_vector( NUMBITS-1 downto 0 ) );
end Decoder;

architecture Behavioral of Decoder is

begin

process(clk)
begin
   if ( clk'event and clk = '1' and read_in = '1' ) then
      if ( rst = '1') then
         output <= "00000000000000000000000000000000";
      else
         case input is
            when "00000" => output <= "00000000000000000000000000000001";
            when "00001" => output <= "00000000000000000000000000000010";
            when "00010" => output <= "00000000000000000000000000000100";
            when "00011" => output <= "00000000000000000000000000001000";
            when "00100" => output <= "00000000000000000000000000010000";
            when "00101" => output <= "00000000000000000000000000100000";
            when "00110" => output <= "00000000000000000000000001000000";
            when "00111" => output <= "00000000000000000000000010000000";
            when "01000" => output <= "00000000000000000000000100000000";
            when "01001" => output <= "00000000000000000000001000000000";
            when "01010" => output <= "00000000000000000000010000000000";
            when "01011" => output <= "00000000000000000000100000000000";
            when "01100" => output <= "00000000000000000001000000000000";
            when "01101" => output <= "00000000000000000010000000000000";
            when "01110" => output <= "00000000000000000100000000000000";
            when "01111" => output <= "00000000000000001000000000000000";
            when "10000" => output <= "00000000000000010000000000000000";
            when "10001" => output <= "00000000000000100000000000000000";
            when "10010" => output <= "00000000000001000000000000000000";
            when "10011" => output <= "00000000000010000000000000000000";
            when "10100" => output <= "00000000000100000000000000000000";
            when "10101" => output <= "00000000001000000000000000000000";
            when "10110" => output <= "00000000010000000000000000000000";
            when "10111" => output <= "00000000100000000000000000000000";
            when "11000" => output <= "00000001000000000000000000000000";
            when "11001" => output <= "00000010000000000000000000000000";
            when "11010" => output <= "00000100000000000000000000000000";
            when "11011" => output <= "00001000000000000000000000000000";
            when "11100" => output <= "00010000000000000000000000000000";
            when "11101" => output <= "00100000000000000000000000000000";
            when "11110" => output <= "01000000000000000000000000000000";
            when "11111" => output <= "10000000000000000000000000000000";
            when others => output <= "00000000000000000000000000000000";
         end case;
      end if;
   end if;
end process;

end Behavioral;

